package enums ;

typedef enum bit [7:0] {  S_0_0,  S_1_0,  S_2_0,  S_3_0,  S_4_0,  S_5_0,  S_6_0,  S_7_0,  S_8_0,  S_9_0,  S_10_0,  S_11_0,  S_12_0,  S_13_0,  S_14_0,  S_15_0,  S_16_0,  S_17_0,  S_18_0,  S_19_0,  S_20_0,  S_21_0,  S_22_0,  S_23_0,  S_24_0,  S_25_0,  S_26_0,  S_27_0,  S_28_0,  S_29_0,  S_30_0,  S_31_0,
                          S_0_1,  S_1_1,  S_2_1,  S_3_1,  S_4_1,  S_5_1,  S_6_1,  S_7_1,  S_8_1,  S_9_1,  S_10_1,  S_11_1,  S_12_1,  S_13_1,  S_14_1,  S_15_1,  S_16_1,  S_17_1,  S_18_1,  S_19_1,  S_20_1,  S_21_1,  S_22_1,  S_23_1,  S_24_1,  S_25_1,  S_26_1,  S_27_1,  S_28_1,  S_29_1,  S_30_1,  S_31_1,
                          S_0_2,  S_1_2,  S_2_2,  S_3_2,  S_4_2,  S_5_2,  S_6_2,  S_7_2,  S_8_2,  S_9_2,  S_10_2,  S_11_2,  S_12_2,  S_13_2,  S_14_2,  S_15_2,  S_16_2,  S_17_2,  S_18_2,  S_19_2,  S_20_2,  S_21_2,  S_22_2,  S_23_2,  S_24_2,  S_25_2,  S_26_2,  S_27_2,  S_28_2,  S_29_2,  S_30_2,  S_31_2,
                          S_0_3,  S_1_3,  S_2_3,  S_3_3,  S_4_3,  S_5_3,  S_6_3,  S_7_3,  S_8_3,  S_9_3,  S_10_3,  S_11_3,  S_12_3,  S_13_3,  S_14_3,  S_15_3,  S_16_3,  S_17_3,  S_18_3,  S_19_3,  S_20_3,  S_21_3,  S_22_3,  S_23_3,  S_24_3,  S_25_3,  S_26_3,  S_27_3,  S_28_3,  S_29_3,  S_30_3,  S_31_3,
                          S_0_4,  S_1_4,  S_2_4,  S_3_4,  S_4_4,  S_5_4,  S_6_4,  S_7_4,  S_8_4,  S_9_4,  S_10_4,  S_11_4,  S_12_4,  S_13_4,  S_14_4,  S_15_4,  S_16_4,  S_17_4,  S_18_4,  S_19_4,  S_20_4,  S_21_4,  S_22_4,  S_23_4,  S_24_4,  S_25_4,  S_26_4,  S_27_4,  S_28_4,  S_29_4,  S_30_4,  S_31_4,
                          S_0_5,  S_1_5,  S_2_5,  S_3_5,  S_4_5,  S_5_5,  S_6_5,  S_7_5,  S_8_5,  S_9_5,  S_10_5,  S_11_5,  S_12_5,  S_13_5,  S_14_5,  S_15_5,  S_16_5,  S_17_5,  S_18_5,  S_19_5,  S_20_5,  S_21_5,  S_22_5,  S_23_5,  S_24_5,  S_25_5,  S_26_5,  S_27_5,  S_28_5,  S_29_5,  S_30_5,  S_31_5,
                          S_0_6,  S_1_6,  S_2_6,  S_3_6,  S_4_6,  S_5_6,  S_6_6,  S_7_6,  S_8_6,  S_9_6,  S_10_6,  S_11_6,  S_12_6,  S_13_6,  S_14_6,  S_15_6,  S_16_6,  S_17_6,  S_18_6,  S_19_6,  S_20_6,  S_21_6,  S_22_6,  S_23_6,  S_24_6,  S_25_6,  S_26_6,  S_27_6,  S_28_6,  S_29_6,  S_30_6,  S_31_6,
                          S_0_7,  S_1_7,  S_2_7,  S_3_7,  S_4_7,  S_5_7,  S_6_7,  S_7_7,  S_8_7,  S_9_7,  S_10_7,  S_11_7,  S_12_7,  S_13_7,  S_14_7,  S_15_7,  S_16_7,  S_17_7,  S_18_7,  S_19_7,  S_20_7,  S_21_7,  S_22_7,  S_23_7,  S_24_7,  S_25_7,  S_26_7,  S_27_7,  S_28_7,  S_29_7,  S_30_7,  S_31_7
                        } data_symbol;

typedef enum bit [7:0] { K_28_0 = 28,
                         K_28_1 = 60,
                         K_28_2 = 92,
                         K_28_3 = 124,
                         K_28_4 = 156,
                         K_28_5 = 188,
                         K_28_6 = 220,
                         K_23_7 = 247,
                         K_27_7 = 251,
                         K_28_7 = 252,
                         K_29_7 = 253,
                         K_30_7 = 254
                        } control_symbol;

endpackage