module assertions_sipo (sipo_if.DUT _if);
    
    //*****************************//
    // TODO: Write Assertions Here //
    //*****************************//

endmodule