package enums ;

typedef enum bit [4:0] {
    S_0_x,  S_1_x,  S_2_x,  S_3_x,  S_4_x,  S_5_x,  S_6_x,  S_7_x,  S_8_x,  S_9_x,  S_10_x,  S_11_x,  S_12_x,  S_13_x,  S_14_x,  S_15_x,  S_16_x,  S_17_x,  S_18_x,  S_19_x,  S_20_x,  S_21_x,  S_22_x,  S_23_x,  S_24_x,  S_25_x,  S_26_x,  S_27_x,  S_28_x,  S_29_x,  S_30_x,  S_31_x
} data_symbol_5;

typedef enum bit [2:0] {
    S_x_0, S_x_1, S_x_2, S_x_3, S_x_4, S_x_5, S_x_6, S_x_7
} data_symbol_3;

typedef enum bit [7:0] {
    S_0_0,  S_1_0,  S_2_0,  S_3_0,  S_4_0,  S_5_0,  S_6_0,  S_7_0,  S_8_0,  S_9_0,  S_10_0,  S_11_0,  S_12_0,  S_13_0,  S_14_0,  S_15_0,  S_16_0,  S_17_0,  S_18_0,  S_19_0,  S_20_0,  S_21_0,  S_22_0,  S_23_0,  S_24_0,  S_25_0,  S_26_0,  S_27_0,  S_28_0,  S_29_0,  S_30_0,  S_31_0,
    S_0_1,  S_1_1,  S_2_1,  S_3_1,  S_4_1,  S_5_1,  S_6_1,  S_7_1,  S_8_1,  S_9_1,  S_10_1,  S_11_1,  S_12_1,  S_13_1,  S_14_1,  S_15_1,  S_16_1,  S_17_1,  S_18_1,  S_19_1,  S_20_1,  S_21_1,  S_22_1,  S_23_1,  S_24_1,  S_25_1,  S_26_1,  S_27_1,  S_28_1,  S_29_1,  S_30_1,  S_31_1,
    S_0_2,  S_1_2,  S_2_2,  S_3_2,  S_4_2,  S_5_2,  S_6_2,  S_7_2,  S_8_2,  S_9_2,  S_10_2,  S_11_2,  S_12_2,  S_13_2,  S_14_2,  S_15_2,  S_16_2,  S_17_2,  S_18_2,  S_19_2,  S_20_2,  S_21_2,  S_22_2,  S_23_2,  S_24_2,  S_25_2,  S_26_2,  S_27_2,  S_28_2,  S_29_2,  S_30_2,  S_31_2,
    S_0_3,  S_1_3,  S_2_3,  S_3_3,  S_4_3,  S_5_3,  S_6_3,  S_7_3,  S_8_3,  S_9_3,  S_10_3,  S_11_3,  S_12_3,  S_13_3,  S_14_3,  S_15_3,  S_16_3,  S_17_3,  S_18_3,  S_19_3,  S_20_3,  S_21_3,  S_22_3,  S_23_3,  S_24_3,  S_25_3,  S_26_3,  S_27_3,  S_28_3,  S_29_3,  S_30_3,  S_31_3,
    S_0_4,  S_1_4,  S_2_4,  S_3_4,  S_4_4,  S_5_4,  S_6_4,  S_7_4,  S_8_4,  S_9_4,  S_10_4,  S_11_4,  S_12_4,  S_13_4,  S_14_4,  S_15_4,  S_16_4,  S_17_4,  S_18_4,  S_19_4,  S_20_4,  S_21_4,  S_22_4,  S_23_4,  S_24_4,  S_25_4,  S_26_4,  S_27_4,  S_28_4,  S_29_4,  S_30_4,  S_31_4,
    S_0_5,  S_1_5,  S_2_5,  S_3_5,  S_4_5,  S_5_5,  S_6_5,  S_7_5,  S_8_5,  S_9_5,  S_10_5,  S_11_5,  S_12_5,  S_13_5,  S_14_5,  S_15_5,  S_16_5,  S_17_5,  S_18_5,  S_19_5,  S_20_5,  S_21_5,  S_22_5,  S_23_5,  S_24_5,  S_25_5,  S_26_5,  S_27_5,  S_28_5,  S_29_5,  S_30_5,  S_31_5,
    S_0_6,  S_1_6,  S_2_6,  S_3_6,  S_4_6,  S_5_6,  S_6_6,  S_7_6,  S_8_6,  S_9_6,  S_10_6,  S_11_6,  S_12_6,  S_13_6,  S_14_6,  S_15_6,  S_16_6,  S_17_6,  S_18_6,  S_19_6,  S_20_6,  S_21_6,  S_22_6,  S_23_6,  S_24_6,  S_25_6,  S_26_6,  S_27_6,  S_28_6,  S_29_6,  S_30_6,  S_31_6,
    S_0_7,  S_1_7,  S_2_7,  S_3_7,  S_4_7,  S_5_7,  S_6_7,  S_7_7,  S_8_7,  S_9_7,  S_10_7,  S_11_7,  S_12_7,  S_13_7,  S_14_7,  S_15_7,  S_16_7,  S_17_7,  S_18_7,  S_19_7,  S_20_7,  S_21_7,  S_22_7,  S_23_7,  S_24_7,  S_25_7,  S_26_7,  S_27_7,  S_28_7,  S_29_7,  S_30_7,  S_31_7
} data_symbol;

typedef enum bit [7:0] {
    K_28_0 = 28,
    K_28_1 = 60,
    K_28_2 = 92,
    K_28_3 = 124,
    K_28_4 = 156,
    K_28_5 = 188,
    K_28_6 = 220,
    K_23_7 = 247,
    K_27_7 = 251,
    K_28_7 = 252,
    K_29_7 = 253,
    K_30_7 = 254
} control_symbol;

typedef enum bit [5:0] {
    E_0_x_p = 6'b000110,
    E_1_x_p = 6'b010001,
    E_2_x_p = 6'b010010,
    E_3_x_p = 6'b100011,
    E_4_x_p = 6'b010100,
    E_5_x_p = 6'b100101,
    E_6_x_p = 6'b100110,
    E_7_x_p = 6'b111000,
    E_8_x_p = 6'b011000,
    E_9_x_p = 6'b101001,
    E_10_x_p = 6'b101010,
    E_11_x_p = 6'b001011,
    E_12_x_p = 6'b101100,
    E_13_x_p = 6'b001101,
    E_14_x_p = 6'b001110,
    E_15_x_p = 6'b000101,
    E_16_x_p = 6'b001001,
    E_17_x_p = 6'b110001,
    E_18_x_p = 6'b110010,
    E_19_x_p = 6'b010011,
    E_20_x_p = 6'b110100,
    E_21_x_p = 6'b010101,
    E_22_x_p = 6'b010110,
    E_23_x_p = 6'b101000,
    E_24_x_p = 6'b001100,
    E_25_x_p = 6'b011001,
    E_26_x_p = 6'b011010,
    E_27_x_p = 6'b100100,
    E_28_x_p = 6'b011100,
    E_29_x_p = 6'b100010,
    E_30_x_p = 6'b100001,
    E_31_x_p = 6'b001010,
    K_28_x_p = 6'b000011
} encoded_word_6_p;

typedef enum bit [5:0] {
    E_0_x_n = 6'b111001,
    E_1_x_n = 6'b101110,
    E_2_x_n = 6'b101101,
    E_3_x_n = 6'b100011,
    E_4_x_n = 6'b101011,
    E_5_x_n = 6'b100101,
    E_6_x_n = 6'b100110,
    E_7_x_n = 6'b000111,
    E_8_x_n = 6'b100111,
    E_9_x_n = 6'b101001,
    E_10_x_n = 6'b101010,
    E_11_x_n = 6'b001011,
    E_12_x_n = 6'b101100,
    E_13_x_n = 6'b001101,
    E_14_x_n = 6'b001110,
    E_15_x_n = 6'b111010,
    E_16_x_n = 6'b110110,
    E_17_x_n = 6'b110001,
    E_18_x_n = 6'b110010,
    E_19_x_n = 6'b010011,
    E_20_x_n = 6'b110100,
    E_21_x_n = 6'b010101,
    E_22_x_n = 6'b010110,
    E_23_x_n = 6'b010111,
    E_24_x_n = 6'b110011,
    E_25_x_n = 6'b011001,
    E_26_x_n = 6'b011010,
    E_27_x_n = 6'b011011,
    E_28_x_n = 6'b011100,
    E_29_x_n = 6'b011101,
    E_30_x_n = 6'b011110,
    E_31_x_n = 6'b110101,
    K_28_x_n = 6'b111100
} encoded_word_6_n;

typedef enum bit [3:0] {
    E_x_0_p  = 4'b0010,
    E_x_1_p  = 4'b1001,
    E_x_2_p  = 4'b1010,
    E_x_3_p  = 4'b1100,
    E_x_4_p  = 4'b0100,
    E_x_5_p  = 4'b0101,
    E_x_6_p  = 4'b0110,
    E_x_P7_p = 4'b1000,
    E_x_A7_p = 4'b0001
} encoded_word_4_p;

typedef enum bit [3:0] {
    K_x_0_p  = 4'b0010,
    K_x_1_p  = 4'b1001,
    K_x_2_p  = 4'b1010,
    K_x_3_p  = 4'b1100,
    K_x_4_p  = 4'b0100,
    K_x_5_p  = 4'b0101,
    K_x_6_p  = 4'b0110,
    K_x_7_p  = 4'b0001
} encoded_control_4_p;

typedef enum bit [3:0] {
    E_x_0_n = 4'b1101,
    E_x_1_n = 4'b1001,
    E_x_2_n = 4'b1010,
    E_x_3_n = 4'b0011,
    E_x_4_n = 4'b1011,
    E_x_5_n = 4'b0101,
    E_x_6_n = 4'b0110,
    E_x_P7_n = 4'b0111,
    E_x_A7_n = 4'b1110
} encoded_word_4_n;

typedef enum bit [3:0] {
    K_x_0_n = 4'b1101,
    K_x_1_n = 4'b0110,
    K_x_2_n = 4'b0101,
    K_x_3_n = 4'b0011,
    K_x_4_n = 4'b1011,
    K_x_5_n = 4'b1010,
    K_x_6_n = 4'b1001,
    K_x_7_n = 4'b1110
} encoded_control_4_n;

typedef enum bit [9:0] {
    E_0_0_p  = {E_x_0_n, E_0_x_p },
    E_1_0_p  = {E_x_0_n, E_1_x_p },
    E_2_0_p  = {E_x_0_n, E_2_x_p },
    E_3_0_p  = {E_x_0_p, E_3_x_p },
    E_4_0_p  = {E_x_0_n, E_4_x_p },
    E_5_0_p  = {E_x_0_p, E_5_x_p },
    E_6_0_p  = {E_x_0_p, E_6_x_p },
    E_7_0_p  = {E_x_0_p, E_7_x_p },
    E_8_0_p  = {E_x_0_n, E_8_x_p },
    E_9_0_p  = {E_x_0_p, E_9_x_p },
    E_10_0_p = {E_x_0_p, E_10_x_p},
    E_11_0_p = {E_x_0_p, E_11_x_p},
    E_12_0_p = {E_x_0_p, E_12_x_p},
    E_13_0_p = {E_x_0_p, E_13_x_p},
    E_14_0_p = {E_x_0_p, E_14_x_p},
    E_15_0_p = {E_x_0_n, E_15_x_p},
    E_16_0_p = {E_x_0_n, E_16_x_p},
    E_17_0_p = {E_x_0_p, E_17_x_p},
    E_18_0_p = {E_x_0_p, E_18_x_p},
    E_19_0_p = {E_x_0_p, E_19_x_p},
    E_20_0_p = {E_x_0_p, E_20_x_p},
    E_21_0_p = {E_x_0_p, E_21_x_p},
    E_22_0_p = {E_x_0_p, E_22_x_p},
    E_23_0_p = {E_x_0_n, E_23_x_p},
    E_24_0_p = {E_x_0_n, E_24_x_p},
    E_25_0_p = {E_x_0_p, E_25_x_p},
    E_26_0_p = {E_x_0_p, E_26_x_p},
    E_27_0_p = {E_x_0_n, E_27_x_p},
    E_28_0_p = {E_x_0_p, E_28_x_p},
    E_29_0_p = {E_x_0_n, E_29_x_p},
    E_30_0_p = {E_x_0_n, E_30_x_p},
    E_31_0_p = {E_x_0_n, E_31_x_p},
    E_0_1_p  = {E_x_1_n, E_0_x_p },
    E_1_1_p  = {E_x_1_n, E_1_x_p },
    E_2_1_p  = {E_x_1_n, E_2_x_p },
    E_3_1_p  = {E_x_1_p, E_3_x_p },
    E_4_1_p  = {E_x_1_n, E_4_x_p },
    E_5_1_p  = {E_x_1_p, E_5_x_p },
    E_6_1_p  = {E_x_1_p, E_6_x_p },
    E_7_1_p  = {E_x_1_p, E_7_x_p },
    E_8_1_p  = {E_x_1_n, E_8_x_p },
    E_9_1_p  = {E_x_1_p, E_9_x_p },
    E_10_1_p = {E_x_1_p, E_10_x_p},
    E_11_1_p = {E_x_1_p, E_11_x_p},
    E_12_1_p = {E_x_1_p, E_12_x_p},
    E_13_1_p = {E_x_1_p, E_13_x_p},
    E_14_1_p = {E_x_1_p, E_14_x_p},
    E_15_1_p = {E_x_1_n, E_15_x_p},
    E_16_1_p = {E_x_1_n, E_16_x_p},
    E_17_1_p = {E_x_1_p, E_17_x_p},
    E_18_1_p = {E_x_1_p, E_18_x_p},
    E_19_1_p = {E_x_1_p, E_19_x_p},
    E_20_1_p = {E_x_1_p, E_20_x_p},
    E_21_1_p = {E_x_1_p, E_21_x_p},
    E_22_1_p = {E_x_1_p, E_22_x_p},
    E_23_1_p = {E_x_1_n, E_23_x_p},
    E_24_1_p = {E_x_1_n, E_24_x_p},
    E_25_1_p = {E_x_1_p, E_25_x_p},
    E_26_1_p = {E_x_1_p, E_26_x_p},
    E_27_1_p = {E_x_1_n, E_27_x_p},
    E_28_1_p = {E_x_1_p, E_28_x_p},
    E_29_1_p = {E_x_1_n, E_29_x_p},
    E_30_1_p = {E_x_1_n, E_30_x_p},
    E_31_1_p = {E_x_1_n, E_31_x_p},
    E_0_2_p  = {E_x_2_n, E_0_x_p },
    E_1_2_p  = {E_x_2_n, E_1_x_p },
    E_2_2_p  = {E_x_2_n, E_2_x_p },
    E_3_2_p  = {E_x_2_p, E_3_x_p },
    E_4_2_p  = {E_x_2_n, E_4_x_p },
    E_5_2_p  = {E_x_2_p, E_5_x_p },
    E_6_2_p  = {E_x_2_p, E_6_x_p },
    E_7_2_p  = {E_x_2_p, E_7_x_p },
    E_8_2_p  = {E_x_2_n, E_8_x_p },
    E_9_2_p  = {E_x_2_p, E_9_x_p },
    E_10_2_p = {E_x_2_p, E_10_x_p},
    E_11_2_p = {E_x_2_p, E_11_x_p},
    E_12_2_p = {E_x_2_p, E_12_x_p},
    E_13_2_p = {E_x_2_p, E_13_x_p},
    E_14_2_p = {E_x_2_p, E_14_x_p},
    E_15_2_p = {E_x_2_n, E_15_x_p},
    E_16_2_p = {E_x_2_n, E_16_x_p},
    E_17_2_p = {E_x_2_p, E_17_x_p},
    E_18_2_p = {E_x_2_p, E_18_x_p},
    E_19_2_p = {E_x_2_p, E_19_x_p},
    E_20_2_p = {E_x_2_p, E_20_x_p},
    E_21_2_p = {E_x_2_p, E_21_x_p},
    E_22_2_p = {E_x_2_p, E_22_x_p},
    E_23_2_p = {E_x_2_n, E_23_x_p},
    E_24_2_p = {E_x_2_n, E_24_x_p},
    E_25_2_p = {E_x_2_p, E_25_x_p},
    E_26_2_p = {E_x_2_p, E_26_x_p},
    E_27_2_p = {E_x_2_n, E_27_x_p},
    E_28_2_p = {E_x_2_p, E_28_x_p},
    E_29_2_p = {E_x_2_n, E_29_x_p},
    E_30_2_p = {E_x_2_n, E_30_x_p},
    E_31_2_p = {E_x_2_n, E_31_x_p},
    E_0_3_p  = {E_x_3_n, E_0_x_p },
    E_1_3_p  = {E_x_3_n, E_1_x_p },
    E_2_3_p  = {E_x_3_n, E_2_x_p },
    E_3_3_p  = {E_x_3_p, E_3_x_p },
    E_4_3_p  = {E_x_3_n, E_4_x_p },
    E_5_3_p  = {E_x_3_p, E_5_x_p },
    E_6_3_p  = {E_x_3_p, E_6_x_p },
    E_7_3_p  = {E_x_3_p, E_7_x_p },
    E_8_3_p  = {E_x_3_n, E_8_x_p },
    E_9_3_p  = {E_x_3_p, E_9_x_p },
    E_10_3_p = {E_x_3_p, E_10_x_p},
    E_11_3_p = {E_x_3_p, E_11_x_p},
    E_12_3_p = {E_x_3_p, E_12_x_p},
    E_13_3_p = {E_x_3_p, E_13_x_p},
    E_14_3_p = {E_x_3_p, E_14_x_p},
    E_15_3_p = {E_x_3_n, E_15_x_p},
    E_16_3_p = {E_x_3_n, E_16_x_p},
    E_17_3_p = {E_x_3_p, E_17_x_p},
    E_18_3_p = {E_x_3_p, E_18_x_p},
    E_19_3_p = {E_x_3_p, E_19_x_p},
    E_20_3_p = {E_x_3_p, E_20_x_p},
    E_21_3_p = {E_x_3_p, E_21_x_p},
    E_22_3_p = {E_x_3_p, E_22_x_p},
    E_23_3_p = {E_x_3_n, E_23_x_p},
    E_24_3_p = {E_x_3_n, E_24_x_p},
    E_25_3_p = {E_x_3_p, E_25_x_p},
    E_26_3_p = {E_x_3_p, E_26_x_p},
    E_27_3_p = {E_x_3_n, E_27_x_p},
    E_28_3_p = {E_x_3_p, E_28_x_p},
    E_29_3_p = {E_x_3_n, E_29_x_p},
    E_30_3_p = {E_x_3_n, E_30_x_p},
    E_31_3_p = {E_x_3_n, E_31_x_p},
    E_0_4_p  = {E_x_4_n, E_0_x_p },
    E_1_4_p  = {E_x_4_n, E_1_x_p },
    E_2_4_p  = {E_x_4_n, E_2_x_p },
    E_3_4_p  = {E_x_4_p, E_3_x_p },
    E_4_4_p  = {E_x_4_n, E_4_x_p },
    E_5_4_p  = {E_x_4_p, E_5_x_p },
    E_6_4_p  = {E_x_4_p, E_6_x_p },
    E_7_4_p  = {E_x_4_p, E_7_x_p },
    E_8_4_p  = {E_x_4_n, E_8_x_p },
    E_9_4_p  = {E_x_4_p, E_9_x_p },
    E_10_4_p = {E_x_4_p, E_10_x_p},
    E_11_4_p = {E_x_4_p, E_11_x_p},
    E_12_4_p = {E_x_4_p, E_12_x_p},
    E_13_4_p = {E_x_4_p, E_13_x_p},
    E_14_4_p = {E_x_4_p, E_14_x_p},
    E_15_4_p = {E_x_4_n, E_15_x_p},
    E_16_4_p = {E_x_4_n, E_16_x_p},
    E_17_4_p = {E_x_4_p, E_17_x_p},
    E_18_4_p = {E_x_4_p, E_18_x_p},
    E_19_4_p = {E_x_4_p, E_19_x_p},
    E_20_4_p = {E_x_4_p, E_20_x_p},
    E_21_4_p = {E_x_4_p, E_21_x_p},
    E_22_4_p = {E_x_4_p, E_22_x_p},
    E_23_4_p = {E_x_4_n, E_23_x_p},
    E_24_4_p = {E_x_4_n, E_24_x_p},
    E_25_4_p = {E_x_4_p, E_25_x_p},
    E_26_4_p = {E_x_4_p, E_26_x_p},
    E_27_4_p = {E_x_4_n, E_27_x_p},
    E_28_4_p = {E_x_4_p, E_28_x_p},
    E_29_4_p = {E_x_4_n, E_29_x_p},
    E_30_4_p = {E_x_4_n, E_30_x_p},
    E_31_4_p = {E_x_4_n, E_31_x_p},
    E_0_5_p  = {E_x_5_n, E_0_x_p },
    E_1_5_p  = {E_x_5_n, E_1_x_p },
    E_2_5_p  = {E_x_5_n, E_2_x_p },
    E_3_5_p  = {E_x_5_p, E_3_x_p },
    E_4_5_p  = {E_x_5_n, E_4_x_p },
    E_5_5_p  = {E_x_5_p, E_5_x_p },
    E_6_5_p  = {E_x_5_p, E_6_x_p },
    E_7_5_p  = {E_x_5_p, E_7_x_p },
    E_8_5_p  = {E_x_5_n, E_8_x_p },
    E_9_5_p  = {E_x_5_p, E_9_x_p },
    E_10_5_p = {E_x_5_p, E_10_x_p},
    E_11_5_p = {E_x_5_p, E_11_x_p},
    E_12_5_p = {E_x_5_p, E_12_x_p},
    E_13_5_p = {E_x_5_p, E_13_x_p},
    E_14_5_p = {E_x_5_p, E_14_x_p},
    E_15_5_p = {E_x_5_n, E_15_x_p},
    E_16_5_p = {E_x_5_n, E_16_x_p},
    E_17_5_p = {E_x_5_p, E_17_x_p},
    E_18_5_p = {E_x_5_p, E_18_x_p},
    E_19_5_p = {E_x_5_p, E_19_x_p},
    E_20_5_p = {E_x_5_p, E_20_x_p},
    E_21_5_p = {E_x_5_p, E_21_x_p},
    E_22_5_p = {E_x_5_p, E_22_x_p},
    E_23_5_p = {E_x_5_n, E_23_x_p},
    E_24_5_p = {E_x_5_n, E_24_x_p},
    E_25_5_p = {E_x_5_p, E_25_x_p},
    E_26_5_p = {E_x_5_p, E_26_x_p},
    E_27_5_p = {E_x_5_n, E_27_x_p},
    E_28_5_p = {E_x_5_p, E_28_x_p},
    E_29_5_p = {E_x_5_n, E_29_x_p},
    E_30_5_p = {E_x_5_n, E_30_x_p},
    E_31_5_p = {E_x_5_n, E_31_x_p},
    E_0_6_p  = {E_x_6_n, E_0_x_p },
    E_1_6_p  = {E_x_6_n, E_1_x_p },
    E_2_6_p  = {E_x_6_n, E_2_x_p },
    E_3_6_p  = {E_x_6_p, E_3_x_p },
    E_4_6_p  = {E_x_6_n, E_4_x_p },
    E_5_6_p  = {E_x_6_p, E_5_x_p },
    E_6_6_p  = {E_x_6_p, E_6_x_p },
    E_7_6_p  = {E_x_6_p, E_7_x_p },
    E_8_6_p  = {E_x_6_n, E_8_x_p },
    E_9_6_p  = {E_x_6_p, E_9_x_p },
    E_10_6_p = {E_x_6_p, E_10_x_p},
    E_11_6_p = {E_x_6_p, E_11_x_p},
    E_12_6_p = {E_x_6_p, E_12_x_p},
    E_13_6_p = {E_x_6_p, E_13_x_p},
    E_14_6_p = {E_x_6_p, E_14_x_p},
    E_15_6_p = {E_x_6_n, E_15_x_p},
    E_16_6_p = {E_x_6_n, E_16_x_p},
    E_17_6_p = {E_x_6_p, E_17_x_p},
    E_18_6_p = {E_x_6_p, E_18_x_p},
    E_19_6_p = {E_x_6_p, E_19_x_p},
    E_20_6_p = {E_x_6_p, E_20_x_p},
    E_21_6_p = {E_x_6_p, E_21_x_p},
    E_22_6_p = {E_x_6_p, E_22_x_p},
    E_23_6_p = {E_x_6_n, E_23_x_p},
    E_24_6_p = {E_x_6_n, E_24_x_p},
    E_25_6_p = {E_x_6_p, E_25_x_p},
    E_26_6_p = {E_x_6_p, E_26_x_p},
    E_27_6_p = {E_x_6_n, E_27_x_p},
    E_28_6_p = {E_x_6_p, E_28_x_p},
    E_29_6_p = {E_x_6_n, E_29_x_p},
    E_30_6_p = {E_x_6_n, E_30_x_p},
    E_31_6_p = {E_x_6_n, E_31_x_p},
    E_0_7_p  = {E_x_P7_n, E_0_x_p },
    E_1_7_p  = {E_x_P7_n, E_1_x_p },
    E_2_7_p  = {E_x_P7_n, E_2_x_p },
    E_3_7_p  = {E_x_P7_p, E_3_x_p },
    E_4_7_p  = {E_x_P7_n, E_4_x_p },
    E_5_7_p  = {E_x_P7_p, E_5_x_p },
    E_6_7_p  = {E_x_P7_p, E_6_x_p },
    E_7_7_p  = {E_x_P7_p, E_7_x_p },
    E_8_7_p  = {E_x_P7_n, E_8_x_p },
    E_9_7_p  = {E_x_P7_p, E_9_x_p },
    E_10_7_p = {E_x_P7_p, E_10_x_p},
    E_11_7_p = {E_x_A7_p, E_11_x_p},
    E_12_7_p = {E_x_P7_p, E_12_x_p},
    E_13_7_p = {E_x_A7_p, E_13_x_p},
    E_14_7_p = {E_x_A7_p, E_14_x_p},
    E_15_7_p = {E_x_P7_n, E_15_x_p},
    E_16_7_p = {E_x_P7_n, E_16_x_p},
    E_17_7_p = {E_x_P7_p, E_17_x_p},
    E_18_7_p = {E_x_P7_p, E_18_x_p},
    E_19_7_p = {E_x_P7_p, E_19_x_p},
    E_20_7_p = {E_x_P7_p, E_20_x_p},
    E_21_7_p = {E_x_P7_p, E_21_x_p},
    E_22_7_p = {E_x_P7_p, E_22_x_p},
    E_23_7_p = {E_x_P7_n, E_23_x_p},
    E_24_7_p = {E_x_P7_n, E_24_x_p},
    E_25_7_p = {E_x_P7_p, E_25_x_p},
    E_26_7_p = {E_x_P7_p, E_26_x_p},
    E_27_7_p = {E_x_P7_n, E_27_x_p},
    E_28_7_p = {E_x_P7_p, E_28_x_p},
    E_29_7_p = {E_x_P7_n, E_29_x_p},
    E_30_7_p = {E_x_P7_n, E_30_x_p},
    E_31_7_p = {E_x_P7_n, E_31_x_p}
} encoded_data_p;

typedef enum bit [9:0] {
    E_0_0_n  = {E_x_0_p, E_0_x_n },
    E_1_0_n  = {E_x_0_p, E_1_x_n },
    E_2_0_n  = {E_x_0_p, E_2_x_n },
    E_3_0_n  = {E_x_0_n, E_3_x_n },
    E_4_0_n  = {E_x_0_p, E_4_x_n },
    E_5_0_n  = {E_x_0_n, E_5_x_n },
    E_6_0_n  = {E_x_0_n, E_6_x_n },
    E_7_0_n  = {E_x_0_n, E_7_x_n },
    E_8_0_n  = {E_x_0_p, E_8_x_n },
    E_9_0_n  = {E_x_0_n, E_9_x_n },
    E_10_0_n = {E_x_0_n, E_10_x_n},
    E_11_0_n = {E_x_0_n, E_11_x_n},
    E_12_0_n = {E_x_0_n, E_12_x_n},
    E_13_0_n = {E_x_0_n, E_13_x_n},
    E_14_0_n = {E_x_0_n, E_14_x_n},
    E_15_0_n = {E_x_0_p, E_15_x_n},
    E_16_0_n = {E_x_0_p, E_16_x_n},
    E_17_0_n = {E_x_0_n, E_17_x_n},
    E_18_0_n = {E_x_0_n, E_18_x_n},
    E_19_0_n = {E_x_0_n, E_19_x_n},
    E_20_0_n = {E_x_0_n, E_20_x_n},
    E_21_0_n = {E_x_0_n, E_21_x_n},
    E_22_0_n = {E_x_0_n, E_22_x_n},
    E_23_0_n = {E_x_0_p, E_23_x_n},
    E_24_0_n = {E_x_0_p, E_24_x_n},
    E_25_0_n = {E_x_0_n, E_25_x_n},
    E_26_0_n = {E_x_0_n, E_26_x_n},
    E_27_0_n = {E_x_0_p, E_27_x_n},
    E_28_0_n = {E_x_0_n, E_28_x_n},
    E_29_0_n = {E_x_0_p, E_29_x_n},
    E_30_0_n = {E_x_0_p, E_30_x_n},
    E_31_0_n = {E_x_0_p, E_31_x_n},
    E_0_1_n  = {E_x_1_p, E_0_x_n },
    E_1_1_n  = {E_x_1_p, E_1_x_n },
    E_2_1_n  = {E_x_1_p, E_2_x_n },
    E_3_1_n  = {E_x_1_n, E_3_x_n },
    E_4_1_n  = {E_x_1_p, E_4_x_n },
    E_5_1_n  = {E_x_1_n, E_5_x_n },
    E_6_1_n  = {E_x_1_n, E_6_x_n },
    E_7_1_n  = {E_x_1_n, E_7_x_n },
    E_8_1_n  = {E_x_1_p, E_8_x_n },
    E_9_1_n  = {E_x_1_n, E_9_x_n },
    E_10_1_n = {E_x_1_n, E_10_x_n},
    E_11_1_n = {E_x_1_n, E_11_x_n},
    E_12_1_n = {E_x_1_n, E_12_x_n},
    E_13_1_n = {E_x_1_n, E_13_x_n},
    E_14_1_n = {E_x_1_n, E_14_x_n},
    E_15_1_n = {E_x_1_p, E_15_x_n},
    E_16_1_n = {E_x_1_p, E_16_x_n},
    E_17_1_n = {E_x_1_n, E_17_x_n},
    E_18_1_n = {E_x_1_n, E_18_x_n},
    E_19_1_n = {E_x_1_n, E_19_x_n},
    E_20_1_n = {E_x_1_n, E_20_x_n},
    E_21_1_n = {E_x_1_n, E_21_x_n},
    E_22_1_n = {E_x_1_n, E_22_x_n},
    E_23_1_n = {E_x_1_p, E_23_x_n},
    E_24_1_n = {E_x_1_p, E_24_x_n},
    E_25_1_n = {E_x_1_n, E_25_x_n},
    E_26_1_n = {E_x_1_n, E_26_x_n},
    E_27_1_n = {E_x_1_p, E_27_x_n},
    E_28_1_n = {E_x_1_n, E_28_x_n},
    E_29_1_n = {E_x_1_p, E_29_x_n},
    E_30_1_n = {E_x_1_p, E_30_x_n},
    E_31_1_n = {E_x_1_p, E_31_x_n},
    E_0_2_n  = {E_x_2_p, E_0_x_n },
    E_1_2_n  = {E_x_2_p, E_1_x_n },
    E_2_2_n  = {E_x_2_p, E_2_x_n },
    E_3_2_n  = {E_x_2_n, E_3_x_n },
    E_4_2_n  = {E_x_2_p, E_4_x_n },
    E_5_2_n  = {E_x_2_n, E_5_x_n },
    E_6_2_n  = {E_x_2_n, E_6_x_n },
    E_7_2_n  = {E_x_2_n, E_7_x_n },
    E_8_2_n  = {E_x_2_p, E_8_x_n },
    E_9_2_n  = {E_x_2_n, E_9_x_n },
    E_10_2_n = {E_x_2_n, E_10_x_n},
    E_11_2_n = {E_x_2_n, E_11_x_n},
    E_12_2_n = {E_x_2_n, E_12_x_n},
    E_13_2_n = {E_x_2_n, E_13_x_n},
    E_14_2_n = {E_x_2_n, E_14_x_n},
    E_15_2_n = {E_x_2_p, E_15_x_n},
    E_16_2_n = {E_x_2_p, E_16_x_n},
    E_17_2_n = {E_x_2_n, E_17_x_n},
    E_18_2_n = {E_x_2_n, E_18_x_n},
    E_19_2_n = {E_x_2_n, E_19_x_n},
    E_20_2_n = {E_x_2_n, E_20_x_n},
    E_21_2_n = {E_x_2_n, E_21_x_n},
    E_22_2_n = {E_x_2_n, E_22_x_n},
    E_23_2_n = {E_x_2_p, E_23_x_n},
    E_24_2_n = {E_x_2_p, E_24_x_n},
    E_25_2_n = {E_x_2_n, E_25_x_n},
    E_26_2_n = {E_x_2_n, E_26_x_n},
    E_27_2_n = {E_x_2_p, E_27_x_n},
    E_28_2_n = {E_x_2_n, E_28_x_n},
    E_29_2_n = {E_x_2_p, E_29_x_n},
    E_30_2_n = {E_x_2_p, E_30_x_n},
    E_31_2_n = {E_x_2_p, E_31_x_n},
    E_0_3_n  = {E_x_3_p, E_0_x_n },
    E_1_3_n  = {E_x_3_p, E_1_x_n },
    E_2_3_n  = {E_x_3_p, E_2_x_n },
    E_3_3_n  = {E_x_3_n, E_3_x_n },
    E_4_3_n  = {E_x_3_p, E_4_x_n },
    E_5_3_n  = {E_x_3_n, E_5_x_n },
    E_6_3_n  = {E_x_3_n, E_6_x_n },
    E_7_3_n  = {E_x_3_n, E_7_x_n },
    E_8_3_n  = {E_x_3_p, E_8_x_n },
    E_9_3_n  = {E_x_3_n, E_9_x_n },
    E_10_3_n = {E_x_3_n, E_10_x_n},
    E_11_3_n = {E_x_3_n, E_11_x_n},
    E_12_3_n = {E_x_3_n, E_12_x_n},
    E_13_3_n = {E_x_3_n, E_13_x_n},
    E_14_3_n = {E_x_3_n, E_14_x_n},
    E_15_3_n = {E_x_3_p, E_15_x_n},
    E_16_3_n = {E_x_3_p, E_16_x_n},
    E_17_3_n = {E_x_3_n, E_17_x_n},
    E_18_3_n = {E_x_3_n, E_18_x_n},
    E_19_3_n = {E_x_3_n, E_19_x_n},
    E_20_3_n = {E_x_3_n, E_20_x_n},
    E_21_3_n = {E_x_3_n, E_21_x_n},
    E_22_3_n = {E_x_3_n, E_22_x_n},
    E_23_3_n = {E_x_3_p, E_23_x_n},
    E_24_3_n = {E_x_3_p, E_24_x_n},
    E_25_3_n = {E_x_3_n, E_25_x_n},
    E_26_3_n = {E_x_3_n, E_26_x_n},
    E_27_3_n = {E_x_3_p, E_27_x_n},
    E_28_3_n = {E_x_3_n, E_28_x_n},
    E_29_3_n = {E_x_3_p, E_29_x_n},
    E_30_3_n = {E_x_3_p, E_30_x_n},
    E_31_3_n = {E_x_3_p, E_31_x_n},
    E_0_4_n  = {E_x_4_p, E_0_x_n },
    E_1_4_n  = {E_x_4_p, E_1_x_n },
    E_2_4_n  = {E_x_4_p, E_2_x_n },
    E_3_4_n  = {E_x_4_n, E_3_x_n },
    E_4_4_n  = {E_x_4_p, E_4_x_n },
    E_5_4_n  = {E_x_4_n, E_5_x_n },
    E_6_4_n  = {E_x_4_n, E_6_x_n },
    E_7_4_n  = {E_x_4_n, E_7_x_n },
    E_8_4_n  = {E_x_4_p, E_8_x_n },
    E_9_4_n  = {E_x_4_n, E_9_x_n },
    E_10_4_n = {E_x_4_n, E_10_x_n},
    E_11_4_n = {E_x_4_n, E_11_x_n},
    E_12_4_n = {E_x_4_n, E_12_x_n},
    E_13_4_n = {E_x_4_n, E_13_x_n},
    E_14_4_n = {E_x_4_n, E_14_x_n},
    E_15_4_n = {E_x_4_p, E_15_x_n},
    E_16_4_n = {E_x_4_p, E_16_x_n},
    E_17_4_n = {E_x_4_n, E_17_x_n},
    E_18_4_n = {E_x_4_n, E_18_x_n},
    E_19_4_n = {E_x_4_n, E_19_x_n},
    E_20_4_n = {E_x_4_n, E_20_x_n},
    E_21_4_n = {E_x_4_n, E_21_x_n},
    E_22_4_n = {E_x_4_n, E_22_x_n},
    E_23_4_n = {E_x_4_p, E_23_x_n},
    E_24_4_n = {E_x_4_p, E_24_x_n},
    E_25_4_n = {E_x_4_n, E_25_x_n},
    E_26_4_n = {E_x_4_n, E_26_x_n},
    E_27_4_n = {E_x_4_p, E_27_x_n},
    E_28_4_n = {E_x_4_n, E_28_x_n},
    E_29_4_n = {E_x_4_p, E_29_x_n},
    E_30_4_n = {E_x_4_p, E_30_x_n},
    E_31_4_n = {E_x_4_p, E_31_x_n},
    E_0_5_n  = {E_x_5_p, E_0_x_n },
    E_1_5_n  = {E_x_5_p, E_1_x_n },
    E_2_5_n  = {E_x_5_p, E_2_x_n },
    E_3_5_n  = {E_x_5_n, E_3_x_n },
    E_4_5_n  = {E_x_5_p, E_4_x_n },
    E_5_5_n  = {E_x_5_n, E_5_x_n },
    E_6_5_n  = {E_x_5_n, E_6_x_n },
    E_7_5_n  = {E_x_5_n, E_7_x_n },
    E_8_5_n  = {E_x_5_p, E_8_x_n },
    E_9_5_n  = {E_x_5_n, E_9_x_n },
    E_10_5_n = {E_x_5_n, E_10_x_n},
    E_11_5_n = {E_x_5_n, E_11_x_n},
    E_12_5_n = {E_x_5_n, E_12_x_n},
    E_13_5_n = {E_x_5_n, E_13_x_n},
    E_14_5_n = {E_x_5_n, E_14_x_n},
    E_15_5_n = {E_x_5_p, E_15_x_n},
    E_16_5_n = {E_x_5_p, E_16_x_n},
    E_17_5_n = {E_x_5_n, E_17_x_n},
    E_18_5_n = {E_x_5_n, E_18_x_n},
    E_19_5_n = {E_x_5_n, E_19_x_n},
    E_20_5_n = {E_x_5_n, E_20_x_n},
    E_21_5_n = {E_x_5_n, E_21_x_n},
    E_22_5_n = {E_x_5_n, E_22_x_n},
    E_23_5_n = {E_x_5_p, E_23_x_n},
    E_24_5_n = {E_x_5_p, E_24_x_n},
    E_25_5_n = {E_x_5_n, E_25_x_n},
    E_26_5_n = {E_x_5_n, E_26_x_n},
    E_27_5_n = {E_x_5_p, E_27_x_n},
    E_28_5_n = {E_x_5_n, E_28_x_n},
    E_29_5_n = {E_x_5_p, E_29_x_n},
    E_30_5_n = {E_x_5_p, E_30_x_n},
    E_31_5_n = {E_x_5_p, E_31_x_n},
    E_0_6_n  = {E_x_6_p, E_0_x_n },
    E_1_6_n  = {E_x_6_p, E_1_x_n },
    E_2_6_n  = {E_x_6_p, E_2_x_n },
    E_3_6_n  = {E_x_6_n, E_3_x_n },
    E_4_6_n  = {E_x_6_p, E_4_x_n },
    E_5_6_n  = {E_x_6_n, E_5_x_n },
    E_6_6_n  = {E_x_6_n, E_6_x_n },
    E_7_6_n  = {E_x_6_n, E_7_x_n },
    E_8_6_n  = {E_x_6_p, E_8_x_n },
    E_9_6_n  = {E_x_6_n, E_9_x_n },
    E_10_6_n = {E_x_6_n, E_10_x_n},
    E_11_6_n = {E_x_6_n, E_11_x_n},
    E_12_6_n = {E_x_6_n, E_12_x_n},
    E_13_6_n = {E_x_6_n, E_13_x_n},
    E_14_6_n = {E_x_6_n, E_14_x_n},
    E_15_6_n = {E_x_6_p, E_15_x_n},
    E_16_6_n = {E_x_6_p, E_16_x_n},
    E_17_6_n = {E_x_6_n, E_17_x_n},
    E_18_6_n = {E_x_6_n, E_18_x_n},
    E_19_6_n = {E_x_6_n, E_19_x_n},
    E_20_6_n = {E_x_6_n, E_20_x_n},
    E_21_6_n = {E_x_6_n, E_21_x_n},
    E_22_6_n = {E_x_6_n, E_22_x_n},
    E_23_6_n = {E_x_6_p, E_23_x_n},
    E_24_6_n = {E_x_6_p, E_24_x_n},
    E_25_6_n = {E_x_6_n, E_25_x_n},
    E_26_6_n = {E_x_6_n, E_26_x_n},
    E_27_6_n = {E_x_6_p, E_27_x_n},
    E_28_6_n = {E_x_6_n, E_28_x_n},
    E_29_6_n = {E_x_6_p, E_29_x_n},
    E_30_6_n = {E_x_6_p, E_30_x_n},
    E_31_6_n = {E_x_6_p, E_31_x_n},
    E_0_7_n  = {E_x_P7_p, E_0_x_n },
    E_1_7_n  = {E_x_P7_p, E_1_x_n },
    E_2_7_n  = {E_x_P7_p, E_2_x_n },
    E_3_7_n  = {E_x_P7_n, E_3_x_n },
    E_4_7_n  = {E_x_P7_p, E_4_x_n },
    E_5_7_n  = {E_x_P7_n, E_5_x_n },
    E_6_7_n  = {E_x_P7_n, E_6_x_n },
    E_7_7_n  = {E_x_P7_n, E_7_x_n },
    E_8_7_n  = {E_x_P7_p, E_8_x_n },
    E_9_7_n  = {E_x_P7_n, E_9_x_n },
    E_10_7_n = {E_x_P7_n, E_10_x_n},
    E_11_7_n = {E_x_P7_n, E_11_x_n},
    E_12_7_n = {E_x_P7_n, E_12_x_n},
    E_13_7_n = {E_x_P7_n, E_13_x_n},
    E_14_7_n = {E_x_P7_n, E_14_x_n},
    E_15_7_n = {E_x_P7_p, E_15_x_n},
    E_16_7_n = {E_x_P7_p, E_16_x_n},
    E_17_7_n = {E_x_A7_n, E_17_x_n},
    E_18_7_n = {E_x_A7_n, E_18_x_n},
    E_19_7_n = {E_x_P7_n, E_19_x_n},
    E_20_7_n = {E_x_A7_n, E_20_x_n},
    E_21_7_n = {E_x_P7_n, E_21_x_n},
    E_22_7_n = {E_x_P7_n, E_22_x_n},
    E_23_7_n = {E_x_P7_p, E_23_x_n},
    E_24_7_n = {E_x_P7_p, E_24_x_n},
    E_25_7_n = {E_x_P7_n, E_25_x_n},
    E_26_7_n = {E_x_P7_n, E_26_x_n},
    E_27_7_n = {E_x_P7_p, E_27_x_n},
    E_28_7_n = {E_x_P7_n, E_28_x_n},
    E_29_7_n = {E_x_P7_p, E_29_x_n},
    E_30_7_n = {E_x_P7_p, E_30_x_n},
    E_31_7_n = {E_x_P7_p, E_31_x_n}
} encoded_data_n;

typedef enum bit [9:0] {
    K_28_0_p = {K_x_0_n, K_28_x_p},
    K_28_1_p = {K_x_1_n, K_28_x_p},
    K_28_2_p = {K_x_2_n, K_28_x_p},
    K_28_3_p = {K_x_3_n, K_28_x_p},
    K_28_4_p = {K_x_4_n, K_28_x_p},
    K_28_5_p = {K_x_5_n, K_28_x_p},
    K_28_6_p = {K_x_6_n, K_28_x_p},
    K_23_7_p = {K_x_7_n, E_23_x_p},
    K_27_7_p = {K_x_7_n, E_27_x_p},
    K_28_7_p = {K_x_7_n, K_28_x_p},
    K_29_7_p = {K_x_7_n, E_29_x_p},
    K_30_7_p = {K_x_7_n, E_30_x_p}
} encoded_control_p;

typedef enum bit [9:0] {
    K_28_0_n = {K_x_0_p, K_28_x_n},
    K_28_1_n = {K_x_1_p, K_28_x_n},
    K_28_2_n = {K_x_2_p, K_28_x_n},
    K_28_3_n = {K_x_3_p, K_28_x_n},
    K_28_4_n = {K_x_4_p, K_28_x_n},
    K_28_5_n = {K_x_5_p, K_28_x_n},
    K_28_6_n = {K_x_6_p, K_28_x_n},
    K_23_7_n = {K_x_7_p, E_23_x_n},
    K_27_7_n = {K_x_7_p, E_27_x_n},
    K_28_7_n = {K_x_7_p, K_28_x_n},
    K_29_7_n = {K_x_7_p, E_29_x_n},
    K_30_7_n = {K_x_7_p, E_30_x_n}
} encoded_control_n;

endpackage