package enums ;

typedef enum bit [7:0] { D_0_0, D_1_0, D_2_0, D_3_0, D_4_0, D_5_0, D_6_0, D_7_0, D_8_0, D_9_0, D_10_0, D_11_0, D_12_0, D_13_0, D_14_0, D_15_0, D_16_0, D_17_0, D_18_0, D_19_0, D_20_0, D_21_0, D_22_0, D_23_0, D_24_0, D_25_0, D_26_0, D_27_0, D_28_0, D_29_0, D_30_0, D_31_0,
                         D_0_1, D_1_1, D_2_1, D_3_1, D_4_1, D_5_1, D_6_1, D_7_1, D_8_1, D_9_1, D_10_1, D_11_1, D_12_1, D_13_1, D_14_1, D_15_1, D_16_1, D_17_1, D_18_1, D_19_1, D_20_1, D_21_1, D_22_1, D_23_1, D_24_1, D_25_1, D_26_1, D_27_1, D_28_1, D_29_1, D_30_1, D_31_1,
                         D_0_2, D_1_2, D_2_2, D_3_2, D_4_2, D_5_2, D_6_2, D_7_2, D_8_2, D_9_2, D_10_2, D_11_2, D_12_2, D_13_2, D_14_2, D_15_2, D_16_2, D_17_2, D_18_2, D_19_2, D_20_2, D_21_2, D_22_2, D_23_2, D_24_2, D_25_2, D_26_2, D_27_2, D_28_2, D_29_2, D_30_2, D_31_2,
                         D_0_3, D_1_3, D_2_3, D_3_3, D_4_3, D_5_3, D_6_3, D_7_3, D_8_3, D_9_3, D_10_3, D_11_3, D_12_3, D_13_3, D_14_3, D_15_3, D_16_3, D_17_3, D_18_3, D_19_3, D_20_3, D_21_3, D_22_3, D_23_3, D_24_3, D_25_3, D_26_3, D_27_3, D_28_3, D_29_3, D_30_3, D_31_3,
                         D_0_4, D_1_4, D_2_4, D_3_4, D_4_4, D_5_4, D_6_4, D_7_4, D_8_4, D_9_4, D_10_4, D_11_4, D_12_4, D_13_4, D_14_4, D_15_4, D_16_4, D_17_4, D_18_4, D_19_4, D_20_4, D_21_4, D_22_4, D_23_4, D_24_4, D_25_4, D_26_4, D_27_4, D_28_4, D_29_4, D_30_4, D_31_4,
                         D_0_5, D_1_5, D_2_5, D_3_5, D_4_5, D_5_5, D_6_5, D_7_5, D_8_5, D_9_5, D_10_5, D_11_5, D_12_5, D_13_5, D_14_5, D_15_5, D_16_5, D_17_5, D_18_5, D_19_5, D_20_5, D_21_5, D_22_5, D_23_5, D_24_5, D_25_5, D_26_5, D_27_5, D_28_5, D_29_5, D_30_5, D_31_5,
                         D_0_6, D_1_6, D_2_6, D_3_6, D_4_6, D_5_6, D_6_6, D_7_6, D_8_6, D_9_6, D_10_6, D_11_6, D_12_6, D_13_6, D_14_6, D_15_6, D_16_6, D_17_6, D_18_6, D_19_6, D_20_6, D_21_6, D_22_6, D_23_6, D_24_6, D_25_6, D_26_6, D_27_6, D_28_6, D_29_6, D_30_6, D_31_6,
                         D_0_7, D_1_7, D_2_7, D_3_7, D_4_7, D_5_7, D_6_7, D_7_7, D_8_7, D_9_7, D_10_7, D_11_7, D_12_7, D_13_7, D_14_7, D_15_7, D_16_7, D_17_7, D_18_7, D_19_7, D_20_7, D_21_7, D_22_7, D_23_7, D_24_7, D_25_7, D_26_7, D_27_7, D_28_7, D_29_7, D_30_7, D_31_7
                        } data_symbol;

endpackage