module assertions_decoder (decoder_if.DUT _if);
    
    //*****************************//
    // TODO: Write Assertions Here //
    //*****************************//

endmodule