module assertions_piso (piso_if.DUT _if);
    
    //*****************************//
    // TODO: Write Assertions Here //
    //*****************************//

endmodule